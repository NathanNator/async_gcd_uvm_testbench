package lc_agent_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "lc_sequence_item.svh"
  `include "lc_cfg.svh"
  `include "lc_monitor.svh"
  `include "lc_driver.svh"
  `include "lc_agent.svh"
  
endpackage: lc_agent_pkg