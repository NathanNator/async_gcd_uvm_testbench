package gcd_test_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import gcd_env_pkg::*;

  `include "gcd_test_base.svh"
  `include "gcd_test.svh"

endpackage: gcd_test_pkg